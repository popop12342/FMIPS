library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity WriteBuffer is
	port (
	);
end WriteBuffer;

architecture WriteBuffer_Arc of WriteBuffer is

begin
	
end WriteBuffer_Arc;